`timescale 1 ns / 1 ns

module ddma_driver_tb #(MEMORY_BUS_WIDTH, FLIT_WIDTH, ADDRESS)(
  input logic clock,
  input logic reset,
  interface_router_port.ROUTER router_if,
  interface_memory.DUT mem_if,
  interface_ddma.TCD ddma_if
);


integer counter = 0;
always @(posedge clock) begin
  counter <= counter + 1;
end


initial begin

  // ============== PE NUM 0 ============== 
  if (ADDRESS == 0) begin

    #0;  // wait 0 cycles

    // source_node:  0
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 6000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 136250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 232500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 328750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 425000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 617500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 713750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 810000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 906250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1098750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1195000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    4096
    // release_time: 1235125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  0
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1237125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1291250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1387500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1580000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1676250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1772500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1868750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2061250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2157500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2253750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2350000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 1 ============== 
  if (ADDRESS == 1) begin

    #0;  // wait 0 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 138250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 140250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 234500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 236500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 330750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 332750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 427000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 429000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 525250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 529250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 619500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 621500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 715750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 717750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 812000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 814000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 908250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 910250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1006500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1010500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1100750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1102750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1197000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1199000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1293250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1295250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1389500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1391500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1487750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1491750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1582000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1584000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1678250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1680250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1774500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1776500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1870750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1872750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1969000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1973000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2063250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2065250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2159500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2161500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2255750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2257750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2352000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2354000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 10 ============== 
  if (ADDRESS == 10) begin

    #0;  // wait 0 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 0
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 108250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 204500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 300750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 397000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 493250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 589500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 685750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 782000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 878250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 974500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1070750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1167000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1263250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1359500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1455750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1552000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1648250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1744500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1840750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1937000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2033250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2129500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2225750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2322000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 11 ============== 
  if (ADDRESS == 11) begin

    #0;  // wait 0 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 44000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 240625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 242625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 523250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 721875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 723875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1004500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1203125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1207125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1485750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1684375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1686375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1967000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 2165625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2167625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 12 ============== 
  if (ADDRESS == 12) begin

    #0;  // wait 0 cycles

    // source_node:  12
    // target_node:  7
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    8192
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 44000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 240625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 721875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  7
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    8192
    // release_time: 1203125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1207125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1684375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 2165625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 13 ============== 
  if (ADDRESS == 13) begin

    #0;  // wait 0 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 136250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 232500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 328750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 425000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 617500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 713750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 810000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 906250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1098750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1195000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1291250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1387500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1580000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1676250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1772500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1868750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2061250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2157500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2253750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2350000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 14 ============== 
  if (ADDRESS == 14) begin

    #0;  // wait 0 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 4000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 100250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 136250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 196500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 232500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 292750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 328750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 389000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 425000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 485250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 581500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 617500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 677750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 713750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 774000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 810000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 870250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 906250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 966500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1062750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1098750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1159000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1195000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1255250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1291250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1351500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1387500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1447750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1544000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1580000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1640250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1676250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1736500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1772500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1832750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1868750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1929000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2025250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2061250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2121500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2157500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2217750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2253750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2314000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2350000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 15 ============== 
  if (ADDRESS == 15) begin

    #0;  // wait 0 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 0
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 136250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 232500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 328750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 425000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 617500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 713750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 810000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 906250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1098750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1195000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1291250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1387500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1580000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1676250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1772500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1868750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2061250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2157500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2253750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2350000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 2 ============== 
  if (ADDRESS == 2) begin

    #0;  // wait 0 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 4000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 242625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 485250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 723875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 966500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1209125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1447750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1686375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1929000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 2167625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 3 ============== 
  if (ADDRESS == 3) begin

    #0;  // wait 0 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 4 ============== 
  if (ADDRESS == 4) begin

    #0;  // wait 0 cycles

    // source_node:  4
    // target_node:  8
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 0, 'Y': 2}
    // data_size:    16384
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 4096;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16384;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #16384;  // wait 8192 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 5 ============== 
  if (ADDRESS == 5) begin

    #0;  // wait 0 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 4000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 42000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 54000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 150250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 240625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 242625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 246500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 342750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 439000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 523250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 535250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 631500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 721875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 723875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 727750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 824000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 920250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1004500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1016500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1112750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  8
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 0, 'Y': 2}
    // data_size:    8192
    // release_time: 1203125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1207125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1209000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1211125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1305250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1401500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1485750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1497750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1594000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1684375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1686375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1690250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1786500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1882750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1967000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1979000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2075250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 2165625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 512;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2048;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #2048;  // wait 1024 cycles

    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 2167625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2171500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2267750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2364000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 6 ============== 
  if (ADDRESS == 6) begin

    #0;  // wait 0 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 50000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 104250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 146250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 200500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 242500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 296750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 338750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 393000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 435000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 489250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 531250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 585500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 627500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 681750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 723750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 778000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 820000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 874250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 916250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 970500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1012500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1066750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1108750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1163000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1205000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1259250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1301250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1355500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1397500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1451750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1493750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1548000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1590000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1644250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1686250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1740500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1782500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1836750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1878750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1933000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1975000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2029250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2071250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2125500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2167500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2221750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2263750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #32768;  // wait 16384 cycles

    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2318000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2360000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 8192;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 32768;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 7 ============== 
  if (ADDRESS == 7) begin

    #0;  // wait 0 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 40000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  3
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 0}
    // data_size:    8192
    // release_time: 42000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 2048;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8192;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #8192;  // wait 4096 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 240625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 721875
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1203125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1684375
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 2165625
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 3;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 1024;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4096;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #4096;  // wait 2048 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end

  // ============== PE NUM 8 ============== 
  if (ADDRESS == 8) begin

    #0;  // wait 0 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 0
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 96250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 136250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    65536
    // release_time: 176000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 16384;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 65536;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #65536;  // wait 32768 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 192500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 232500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    65536
    // release_time: 272000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 16384;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 65536;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #65536;  // wait 32768 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 288750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 328750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 385000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 425000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 481250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 521250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 577500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 617500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 673750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 713750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 770000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 810000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 866250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 906250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 962500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1002500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1058750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1098750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1155000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1195000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1251250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1291250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1347500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1387500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    65536
    // release_time: 1427125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 16384;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 65536;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #65536;  // wait 32768 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1443750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1483750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    65536
    // release_time: 1523125
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << 16) & 1;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 16384;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 65536;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #65536;  // wait 32768 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1540000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1580000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1636250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1676250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1732500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1772500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1828750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1868750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1925000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1965000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2021250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2061250
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2117500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2157500
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2213750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2253750
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2310000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 0;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
    #153600;  // wait 76800 cycles

    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2350000
    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << 16) & 2;  // header flit
    mem_if.addr_in = 'h0;

    #2;
    mem_if.enable_in = 1;
    mem_if.wb_in = 1;
    mem_if.data_in = 38400;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h4;

    #2;
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 153600;
    ddma_if.cmd_in = 1;

    mem_if.wb_in = 0;  // lock memory write


    #2;
  end



end

endmodule

