module ddma_driver_tb1 #()(
  input logic clock,
  input logic reset,
  interface_router_port.ROUTER router_if,
  interface_memory.DUT mem_if,
  interface_ddma.TCD ddma_if
);


integer counter = 0;
always @(posedge clock) begin
  counter <= counter + 1;
end


initial begin

  router_if.clock_tx = clock;
  router_if.data_o = counter;
  #0;  // wait 0 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 40000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 138250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 140250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 234500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 236500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 330750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 332750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 427000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 429000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 525250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 529250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 619500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 621500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 715750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 717750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 812000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 814000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 908250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 910250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1006500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1010500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1100750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1102750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1197000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1199000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1293250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1295250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1389500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1391500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1487750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1491750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1582000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1584000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1678250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1680250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1774500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1776500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1870750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1872750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 1969000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 1973000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 2063250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 2065250
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 2159500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 2161500
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 2255750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 2257750
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #8192;  // wait 4096 cycles

  // source_node:  1
  // target_node:  5
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 1, 'Y': 1}
  // data_size:    2048
  // release_time: 2352000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (1 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 512;  // 2048 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 2048;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
  #2048;  // wait 1024 cycles

  // source_node:  1
  // target_node:  6
  // source_xy:    {'X': 1, 'Y': 0}
  // target_xy:    {'X': 2, 'Y': 1}
  // data_size:    8192
  // release_time: 2354000
  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = (2 << 16) & 1;  // header flit
  mem_if.addr_in = 'h0;

  #2;
  mem_if.enable_in = 1;
  mem_if.wb_in = 1;
  mem_if.data_in = 2048;  // 8192 bytes, size flit
  mem_if.addr_in = 'h0 + 'h4;

  #2;
  ddma_if.addr_in = 'h0;
  ddma_if.nbytes = 8192;
  ddma_if.cmd_in = 1;

  mem_if.wb_in = 0;  // lock memory write


  #2;
end

endmodule

