`timescale 1ns/10ps

module ddma_driver_tb #(MEMORY_BUS_WIDTH, FLIT_WIDTH, ADDRESS)(
  input logic clock,
  input logic reset,
  interface_memory.DUT mem_if,
  interface_ddma.TCD ddma_if
);


integer counter = 0;
always @(posedge clock) begin
  counter <= counter + 1;
end


initial begin

  // delay to handle initialization offset
  mem_if.enable_in = 1;
  ddma_if.addr_in = 0;
  ddma_if.nbytes_in = 0;
  ddma_if.cmd_in = 0;
  // ============== PE NUM 0 ============== 
  if (ADDRESS == 0) begin

    // pkt name:     f31:0
    // source_node:  0
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 6000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #6098; // skipt to 6000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:0
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #33997; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f1:0
    // source_node:  0
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    4096
    // release_time: 80000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 80000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:1
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:2
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:3
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:4
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:5
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:6
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:7
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:8
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:9
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:10
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:11
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:12
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f1:1
    // source_node:  0
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    4096
    // release_time: 1235125
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40122; // skipt to 1235125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f31:1
    // source_node:  0
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1237125
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1237125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:13
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54122; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:14
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:15
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:16
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:17
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:18
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:19
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:20
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:21
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:22
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:23
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f12:24
    // source_node:  0
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2350000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2350000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 1 ============== 
  if (ADDRESS == 1) begin

    // pkt name:     f20:0
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:1
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 138250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #98247; // skipt to 138250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:1
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 140250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 140250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:2
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 234500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 234500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:2
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 236500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 236500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:3
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 330750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 330750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:3
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 332750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 332750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:4
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 427000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 427000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:4
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 429000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 429000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:5
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 525250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 525250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:5
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 529250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 529250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:6
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 619500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90247; // skipt to 619500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:6
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 621500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 621500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:7
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 715750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 715750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:7
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 717750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 717750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:8
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 812000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 812000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:8
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 814000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 814000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:9
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 908250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 908250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:9
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 910250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 910250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:10
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1006500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1006500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:10
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1010500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1010500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:11
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1100750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90247; // skipt to 1100750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:11
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1102750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1102750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:12
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1197000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1197000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:12
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1199000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1199000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:13
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1293250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1293250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:13
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1295250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1295250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:14
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1389500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1389500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:14
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1391500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1391500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:15
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1487750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1487750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:15
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1491750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1491750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:16
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1582000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90247; // skipt to 1582000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:16
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1584000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1584000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:17
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1678250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1678250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:17
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1680250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1680250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:18
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1774500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1774500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:18
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1776500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1776500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:19
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1870750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 1870750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:19
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1872750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1872750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:20
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1969000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1969000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:20
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1973000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1973000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:21
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2063250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90247; // skipt to 2063250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:21
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2065250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2065250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:22
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2159500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 2159500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:22
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2161500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2161500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:23
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2255750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 2255750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:23
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2257750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2257750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f10:24
    // source_node:  1
    // target_node:  5
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2352000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94247; // skipt to 2352000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f20:24
    // source_node:  1
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2354000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2354000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 10 ============== 
  if (ADDRESS == 10) begin

    // pkt name:     f30:0
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 0
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #98; // skipt to 0
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:1
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:1
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 108250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 108250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:2
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:2
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 204500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 204500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:3
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:3
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 300750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 300750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:4
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:4
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 397000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 397000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:5
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:5
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 493250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 493250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:6
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:6
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 589500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 589500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:7
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:7
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 685750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 685750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:8
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:8
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 782000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 782000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:9
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:9
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 878250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 878250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:10
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:10
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 974500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 974500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:11
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:11
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1070750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1070750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:12
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:12
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1167000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1167000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:13
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:13
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1263250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1263250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:14
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:14
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1359500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1359500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:15
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:15
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1455750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1455750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:16
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:16
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1552000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1552000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:17
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:17
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1648250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1648250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:18
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:18
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1744500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1744500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:19
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:19
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1840750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1840750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:20
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:20
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1937000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1937000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:21
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:21
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2033250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 2033250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:22
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:22
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2129500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 2129500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:23
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:23
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2225750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 2225750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f30:24
    // source_node:  10
    // target_node:  4
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    16384
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #84247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f26:24
    // source_node:  10
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2322000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 2322000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 11 ============== 
  if (ADDRESS == 11) begin

    // pkt name:     f6:0
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:0
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 44000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 44000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:1
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #52247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:2
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:1
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 240625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 240625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:1
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 242625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 242625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:3
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:4
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:5
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:2
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:2
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 523250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 523250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:6
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:7
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:3
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 721875
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 721875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:3
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 723875
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 723875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:8
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:9
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:10
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:4
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:4
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1004500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1004500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:11
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:12
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:5
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1203125
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1203125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:5
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1207125
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1207125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:13
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #44122; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:14
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:15
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:6
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:6
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1485750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1485750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:16
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:17
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:7
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1684375
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1684375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:7
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1686375
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1686375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:18
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:19
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:20
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:8
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:8
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1967000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1967000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:21
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:22
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f37:9
    // source_node:  11
    // target_node:  7
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    4096
    // release_time: 2165625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 2165625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f6:9
    // source_node:  11
    // target_node:  5
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2167625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2167625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:23
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f18:24
    // source_node:  11
    // target_node:  10
    // source_xy:    {'X': 3, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 12 ============== 
  if (ADDRESS == 12) begin

    // pkt name:     f34:0
    // source_node:  12
    // target_node:  7
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    8192
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:0
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 44000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 44000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:1
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #52247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:2
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:1
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 240625
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 240625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:3
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:4
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:5
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:2
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:6
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:7
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:3
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 721875
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 721875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:8
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:9
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:10
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:4
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:11
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:12
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f34:1
    // source_node:  12
    // target_node:  7
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    8192
    // release_time: 1203125
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1203125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:5
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1207125
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1207125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:13
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #44122; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:14
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:15
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:6
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:16
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:17
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:7
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1684375
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1684375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:18
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:19
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:20
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:8
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:21
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:22
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f32:9
    // source_node:  12
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    4096
    // release_time: 2165625
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 2165625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:23
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f15:24
    // source_node:  12
    // target_node:  13
    // source_xy:    {'X': 0, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 13 ============== 
  if (ADDRESS == 13) begin

    // pkt name:     f23:1
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #136348; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:2
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:3
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:4
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:5
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:6
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:7
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:8
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:9
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:10
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:11
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:12
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:13
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:14
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:15
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:16
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:17
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:18
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:19
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:20
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:21
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:22
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:23
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f23:24
    // source_node:  13
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2350000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2350000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 14 ============== 
  if (ADDRESS == 14) begin

    // pkt name:     f27:0
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 4000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #4098; // skipt to 4000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:1
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 100250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 100250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:1
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:2
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 196500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 196500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:2
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:3
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 292750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 292750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:3
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:4
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 389000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 389000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:4
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:5
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 485250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 485250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:5
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:6
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 581500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 581500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:6
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:7
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 677750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 677750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:7
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:8
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 774000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 774000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:8
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:9
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 870250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 870250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:9
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:10
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 966500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 966500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:10
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:11
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1062750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1062750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:11
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:12
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1159000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1159000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:12
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:13
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1255250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1255250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:13
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:14
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1351500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1351500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:14
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:15
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1447750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1447750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:15
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:16
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1544000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1544000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:16
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:17
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1640250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1640250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:17
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:18
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1736500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1736500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:18
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:19
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1832750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1832750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:19
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:20
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1929000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 1929000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:20
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:21
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2025250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 2025250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:21
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:22
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2121500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 2121500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:22
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:23
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2217750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 2217750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:23
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f27:24
    // source_node:  14
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2314000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #60247; // skipt to 2314000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f11:24
    // source_node:  14
    // target_node:  5
    // source_xy:    {'X': 2, 'Y': 3}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    2048
    // release_time: 2350000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #35997; // skipt to 2350000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 15 ============== 
  if (ADDRESS == 15) begin

    // pkt name:     f9:0
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 0
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #98; // skipt to 0
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:1
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:1
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:2
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:2
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:3
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:3
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:4
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:4
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:5
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:5
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:6
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:6
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:7
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:7
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:8
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:8
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:9
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:9
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:10
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:10
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:11
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:11
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:12
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:12
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:13
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:13
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:14
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:14
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:15
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:15
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:16
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:16
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:17
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:17
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:18
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:18
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:19
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:19
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:20
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:20
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:21
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:21
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:22
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:22
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:23
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:23
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f9:24
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f19:24
    // source_node:  15
    // target_node:  14
    // source_xy:    {'X': 3, 'Y': 3}
    // target_xy:    {'X': 2, 'Y': 3}
    // data_size:    153600
    // release_time: 2350000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2350000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 2 ============== 
  if (ADDRESS == 2) begin

    // pkt name:     f35:0
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 4000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #4098; // skipt to 4000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:1
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #92247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:2
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:1
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 242625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #50122; // skipt to 242625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:3
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:4
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:5
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:2
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 485250
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 485250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:6
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #92247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:7
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:3
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 723875
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #50122; // skipt to 723875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:8
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:9
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:10
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:4
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 966500
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 966500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:11
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #92247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:12
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:5
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1209125
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54122; // skipt to 1209125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:13
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #42122; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:14
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:15
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:6
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1447750
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1447750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:16
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #92247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:17
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:7
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1686375
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #50122; // skipt to 1686375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:18
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:19
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:20
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:8
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 1929000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1929000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:21
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #92247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:22
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f35:9
    // source_node:  2
    // target_node:  7
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 3, 'Y': 1}
    // data_size:    2048
    // release_time: 2167625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #50122; // skipt to 2167625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:23
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #46122; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f24:24
    // source_node:  2
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 0}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 3 ============== 
  if (ADDRESS == 3) begin

    // pkt name:     f16:1
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96348; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:2
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:3
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:4
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:5
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:6
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:7
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:8
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:9
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:10
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:11
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:12
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:13
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:14
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:15
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:16
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:17
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:18
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:19
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:20
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:21
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:22
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:23
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f16:24
    // source_node:  3
    // target_node:  2
    // source_xy:    {'X': 3, 'Y': 0}
    // target_xy:    {'X': 2, 'Y': 0}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 4 ============== 
  if (ADDRESS == 4) begin

    // pkt name:     f33:0
    // source_node:  4
    // target_node:  8
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 0, 'Y': 2}
    // data_size:    16384
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 4097;  // 16384 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 4099;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:1
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:2
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:3
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:4
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:5
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:6
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:7
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:8
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:9
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:10
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:11
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:12
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:13
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:14
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:15
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:16
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:17
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:18
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:19
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:20
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:21
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:22
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:23
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f13:24
    // source_node:  4
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 5 ============== 
  if (ADDRESS == 5) begin

    // pkt name:     f5:0
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 4000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #4098; // skipt to 4000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:0
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 42000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #37997; // skipt to 42000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:0
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 54000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 54000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:1
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 150250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 150250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:1
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 240625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90372; // skipt to 240625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:1
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 242625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 242625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:2
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 246500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3872; // skipt to 246500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:3
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 342750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 342750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:4
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 439000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 439000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:2
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #42247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:2
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 523250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 523250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:5
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 535250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 535250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:6
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 631500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 631500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:3
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 721875
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90372; // skipt to 721875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:3
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 723875
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 723875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:7
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 727750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3872; // skipt to 727750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:8
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 824000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 824000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:9
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 920250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 920250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:4
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #42247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:4
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1004500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1004500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:10
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1016500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1016500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:11
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1112750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1112750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f2:1
    // source_node:  5
    // target_node:  8
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 0, 'Y': 2}
    // data_size:    8192
    // release_time: 1203125
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90372; // skipt to 1203125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:5
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1207125
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3997; // skipt to 1207125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:12
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1209000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1872; // skipt to 1209000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:5
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1211125
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #2122; // skipt to 1211125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:13
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1305250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #94122; // skipt to 1305250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:14
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1401500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1401500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:6
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #42247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:6
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1485750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1485750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:15
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1497750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1497750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:16
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1594000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1594000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:7
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1684375
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90372; // skipt to 1684375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:7
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1686375
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 1686375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:17
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1690250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3872; // skipt to 1690250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:18
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1786500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1786500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:19
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1882750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1882750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:8
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #42247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:8
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1967000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1967000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:20
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1979000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #11997; // skipt to 1979000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:21
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2075250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2075250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f5:9
    // source_node:  5
    // target_node:  15
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 3}
    // data_size:    2048
    // release_time: 2165625
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 513;  // 2048 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #90372; // skipt to 2165625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 515;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f7:9
    // source_node:  5
    // target_node:  13
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 2167625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 2167625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:22
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2171500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #3872; // skipt to 2171500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:23
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2267750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2267750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f21:24
    // source_node:  5
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2364000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2364000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 6 ============== 
  if (ADDRESS == 6) begin

    // pkt name:     f28:0
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 50000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #50098; // skipt to 50000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:1
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 104250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 104250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:1
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 146250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 146250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:2
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 200500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 200500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:2
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 242500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 242500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:3
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 296750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 296750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:3
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 338750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 338750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:4
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 393000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 393000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:4
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 435000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 435000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:5
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 489250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 489250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:5
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 531250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 531250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:6
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 585500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 585500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:6
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 627500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 627500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:7
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 681750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 681750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:7
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 723750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 723750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:8
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 778000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 778000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:8
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 820000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 820000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:9
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 874250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 874250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:9
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 916250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 916250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:10
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 970500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 970500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:10
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1012500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1012500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:11
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1066750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1066750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:11
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1108750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1108750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:12
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1163000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1163000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:12
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1205000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1205000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:13
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1259250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1259250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:13
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1301250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1301250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:14
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1355500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1355500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:14
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1397500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1397500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:15
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1451750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1451750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:15
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1493750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1493750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:16
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1548000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1548000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:16
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1590000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1590000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:17
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1644250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1644250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:17
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1686250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1686250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:18
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1740500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1740500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:18
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1782500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1782500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:19
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1836750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1836750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:19
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1878750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1878750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:20
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 1933000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 1933000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:20
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1975000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 1975000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:21
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2029250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 2029250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:21
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2071250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 2071250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:22
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2125500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 2125500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:22
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2167500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 2167500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:23
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2221750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 2221750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:23
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2263750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 2263750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f25:24
    // source_node:  6
    // target_node:  9
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    8192
    // release_time: 2318000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 2318000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f28:24
    // source_node:  6
    // target_node:  10
    // source_xy:    {'X': 2, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2360000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #41997; // skipt to 2360000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 7 ============== 
  if (ADDRESS == 7) begin

    // pkt name:     f38:0
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f36:0
    // source_node:  7
    // target_node:  3
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 3, 'Y': 0}
    // data_size:    8192
    // release_time: 42000
    mem_if.wb_in = 1;
    mem_if.data_in = (3 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #1997; // skipt to 42000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:1
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #54247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:2
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:1
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 240625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 240625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:3
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:4
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:5
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:2
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:6
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:7
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:3
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 721875
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 721875
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:8
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:9
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:10
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:4
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:11
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:12
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:5
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1203125
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1203125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:13
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:14
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:15
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:6
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:16
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:17
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:7
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1684375
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1684375
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:18
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:19
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:20
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:8
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:21
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:22
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f38:9
    // source_node:  7
    // target_node:  13
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 1, 'Y': 3}
    // data_size:    4096
    // release_time: 2165625
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 3;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 1025;  // 4096 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 2165625
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 1027;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:23
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #48122; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f17:24
    // source_node:  7
    // target_node:  6
    // source_xy:    {'X': 3, 'Y': 1}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 8 ============== 
  if (ADDRESS == 8) begin

    // pkt name:     f8:0
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 0
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #98; // skipt to 0
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:1
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 96250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 96250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:1
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f3:0
    // source_node:  8
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    65536
    // release_time: 176000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 16385;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39747; // skipt to 176000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16387;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:2
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 192500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #16497; // skipt to 192500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:2
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f4:0
    // source_node:  8
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    65536
    // release_time: 272000
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 16385;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39497; // skipt to 272000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16387;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:3
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 288750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #16747; // skipt to 288750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:3
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:4
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 385000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 385000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:4
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:5
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 481250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 481250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:5
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:6
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 577500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 577500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:6
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:7
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 673750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 673750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:7
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:8
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 770000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 770000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:8
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:9
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 866250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 866250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:9
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:10
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 962500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 962500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:10
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:11
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1058750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1058750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:11
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:12
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1155000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1155000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:12
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:13
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1251250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1251250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:13
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:14
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1347500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1347500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:14
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f3:1
    // source_node:  8
    // target_node:  5
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 1}
    // data_size:    65536
    // release_time: 1427125
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 16385;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39622; // skipt to 1427125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16387;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:15
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1443750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #16622; // skipt to 1443750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:15
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f4:1
    // source_node:  8
    // target_node:  4
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 0, 'Y': 1}
    // data_size:    65536
    // release_time: 1523125
    mem_if.wb_in = 1;
    mem_if.data_in = (0 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 16385;  // 65536 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39372; // skipt to 1523125
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 16387;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:16
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1540000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #16872; // skipt to 1540000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:16
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:17
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1636250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1636250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:17
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:18
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1732500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1732500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:18
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:19
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1828750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1828750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:19
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:20
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 1925000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 1925000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:20
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:21
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2021250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2021250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:21
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:22
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2117500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2117500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:22
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:23
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2213750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2213750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:23
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f8:24
    // source_node:  8
    // target_node:  1
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 0}
    // data_size:    153600
    // release_time: 2310000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 0;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #56247; // skipt to 2310000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f14:24
    // source_node:  8
    // target_node:  9
    // source_xy:    {'X': 0, 'Y': 2}
    // target_xy:    {'X': 1, 'Y': 2}
    // data_size:    153600
    // release_time: 2350000
    mem_if.wb_in = 1;
    mem_if.data_in = (1 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 38401;  // 153600 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #39997; // skipt to 2350000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 38403;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end

  // ============== PE NUM 9 ============== 
  if (ADDRESS == 9) begin

    // pkt name:     f29:0
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 40000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #40098; // skipt to 40000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:1
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 136250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 136250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:1
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 146250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 146250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:2
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 232500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 232500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:2
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 242500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 242500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:3
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 328750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 328750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:3
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 338750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 338750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:4
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 425000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 425000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:4
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 435000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 435000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:5
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 521250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 521250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:5
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 531250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 531250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:6
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 617500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 617500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:6
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 627500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 627500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:7
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 713750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 713750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:7
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 723750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 723750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:8
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 810000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 810000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:8
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 820000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 820000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:9
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 906250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 906250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:9
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 916250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 916250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:10
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1002500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1002500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:10
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1012500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1012500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:11
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1098750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1098750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:11
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1108750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1108750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:12
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1195000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1195000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:12
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1205000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1205000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:13
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1291250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1291250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:13
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1301250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1301250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:14
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1387500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1387500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:14
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1397500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1397500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:15
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1483750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1483750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:15
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1493750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1493750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:16
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1580000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1580000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:16
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1590000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1590000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:17
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1676250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1676250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:17
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1686250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1686250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:18
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1772500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1772500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:18
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1782500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1782500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:19
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1868750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1868750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:19
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1878750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1878750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:20
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 1965000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 1965000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:20
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 1975000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 1975000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:21
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2061250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 2061250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:21
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2071250
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 2071250
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:22
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2157500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 2157500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:22
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2167500
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 2167500
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f29:23
    // source_node:  9
    // target_node:  10
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 2}
    // data_size:    32768
    // release_time: 2253750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 2;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 8193;  // 32768 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #86247; // skipt to 2253750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 8195;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:23
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2263750
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #9997; // skipt to 2263750
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
    // pkt name:     f22:24
    // source_node:  9
    // target_node:  6
    // source_xy:    {'X': 1, 'Y': 2}
    // target_xy:    {'X': 2, 'Y': 1}
    // data_size:    8192
    // release_time: 2360000
    mem_if.wb_in = 1;
    mem_if.data_in = (2 << (FLIT_WIDTH / 4)) | 1;
    mem_if.addr_in = 'h0;
    #1;

    mem_if.wb_in = 1;
    mem_if.data_in = 2049;  // 8192 bytes, size flit
    mem_if.addr_in = 'h0 + 'h1;
    #1;

    mem_if.wb_in = 0;  // lock memory write


    #96247; // skipt to 2360000
    ddma_if.addr_in = 'h0;
    ddma_if.nbytes_in = 2051;
    ddma_if.cmd_in = 1;
    #1;

    ddma_if.addr_in = 0;
    ddma_if.nbytes_in = 0;
    ddma_if.cmd_in = 0; 
  end



end

endmodule

